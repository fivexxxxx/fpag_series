
/*
"="   阻塞赋值运算符
"<="  非阻塞赋值运算符

阻塞赋值运算符：阻塞赋值运算符在执行赋值操作时，会暂停当前进程的执行，直到赋值完成。
这意味着在当前时间步内，其他进程无法访问或修改被赋值的变量，直到该变量的值更新完毕。

非阻塞赋值运算符：非阻塞赋值运算符在执行赋值操作时，不会暂停当前进程的执行。
这意味着在当前时间步内，其他进程仍然可以访问或修改被赋值的变量，即使该变量的值尚未更新完毕。




*/
`timescale 1ns / 1ps

module tb_ex;
reg                     a               ;
reg                     b               ;   
reg                     c               ;
reg                     d               ;
reg                     e               ;
reg                     f               ;
//阻塞赋值与非阻塞赋值的区别：
//阻塞赋值

initial begin
    a = 0;
    b = 1;
    c = a+b;
end

//非阻塞赋值

initial begin
    d <= 0;
    e <= 1;
    f <= d+e;
end


endmodule